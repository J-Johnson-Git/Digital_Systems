`timescale 1ns / 1ps


module uart_tx_tb
(
    
);
endmodule
